        -- addi $r1 $r0 0xfefe
        0 => x"20",
        1 => x"01",
        2 => x"fe",
        3 => x"fe",

        -- addi $r2 $r0 0xcece
        4 => x"20",
        5 => x"02",
        6 => x"ce",
        7 => x"ce",

        -- nop
        8 => x"00",
        9 => x"00",
        10 => x"00",
        11 => x"00",

        -- nop
        12 => x"00",
        13 => x"00",
        14 => x"00",
        15 => x"00",

        -- sw $r1 16($r0)
        16 => x"ac",
        17 => x"01",
        18 => x"00",
        19 => x"10",

        -- andi $r3 $r2 0x8
        20 => x"30",
        21 => x"43",
        22 => x"00",
        23 => x"08",

        -- ori $r4 $r2 0x7
        24 => x"34",
        25 => x"44",
        26 => x"00",
        27 => x"07",

        -- xori $r5 $r2 0x7
        28 => x"38",
        29 => x"45",
        30 => x"00",
        31 => x"07",

        -- lw $r6 16($r0)
        32 => x"8c",
        33 => x"06",
        34 => x"00",
        35 => x"10",

        -- multu $r7 $r1 $r2
        36 => x"00",
        37 => x"22",
        38 => x"38",
        39 => x"19",

        -- sll $r8 $r1 $r3
        40 => x"00",
        41 => x"23",
        42 => x"40",
        43 => x"00",

        -- sra $r9 $r2 $r3
        44 => x"00",
        45 => x"43",
        46 => x"48",
        47 => x"03",

        -- srl $r10 $r2 $r3
        48 => x"00",
        49 => x"43",
        50 => x"50",
        51 => x"02",

        -- sub $r11 $r1 $r2
        52 => x"00",
        53 => x"22",
        54 => x"58",
        55 => x"22",

        -- add $r12 $r1 $r2
        56 => x"00",
        57 => x"22",
        58 => x"60",
        59 => x"20",

        -- and $r13 $r1 $r2
        60 => x"00",
        61 => x"22",
        62 => x"68",
        63 => x"24",

        -- or $r14 $r1 $r2
        64 => x"00",
        65 => x"22",
        66 => x"70",
        67 => x"25",

        -- xor $r15 $r1 $r2
        68 => x"00",
        69 => x"22",
        70 => x"78",
        71 => x"26",

